module ghost_motion();


endmodule